
/******************************************************************
* Description
*
* Debouncer
*
* Author: Juan Antonio Serrano Gomez
* email : antonio.serrano@cinvestav.mx
* Date  :	09/06/2023
******************************************************************/

module debouncer(input pb_1, clk,output pb_out);
	wire slow_clk_en;
	wire Q1,Q2,Q2_bar,Q0;
	
	clock_enable u1(clk,slow_clk_en);
	my_dff_en d0(clk,slow_clk_en,pb_1,Q0);
	my_dff_en d1(clk,slow_clk_en,Q0,Q1);
	my_dff_en d2(clk,slow_clk_en,Q1,Q2);
	
//	assign Q2_bar = ~;
	assign pb_out = Q2;
endmodule


// Slow clock enable for debouncing button 
module clock_enable(input Clk_100M,output slow_clk_en);
    reg [26:0]counter=0;
    always @(posedge Clk_100M)
    begin
       counter <= (counter>=249999)?0:counter+1;
    end

    assign slow_clk_en = (counter == 249999)?1'b1:1'b0;
endmodule

// D-flip-flop with clock enable signal for debouncing module 
module my_dff_en(input DFF_CLOCK, clock_enable,D, output reg Q=0);
	always @ (posedge DFF_CLOCK) begin
	if(clock_enable==1)	Q <= D;
    end
endmodule 
