

//Demultiplexor 1 a 4
module mux4to1_case (a,sel,y);
	input [3:0] a;
	input [1:0] sel;
	output reg y;
	
	always_comb begin
		case(sel)
		2'b00: begin y = a[0]; end
		2'b01: begin y = a[1]; end
		2'b10: begin y = a[2]; end
		2'b11: begin y = a[3]; end
		default: y = 1'b0;endcase
	end 
endmodule
	