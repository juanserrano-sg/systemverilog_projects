module TBej4_BCDto7;
logic [3:0] a;
logic [6:0] y;

ej4_BCDto7 dut(.a(a), .y(y)); 
	initial begin
		a = 0;
		#100;
		a = 1;
		#100;
		a = 2;
		#100;
		a = 3;
		#100;
		a = 4;
		#100;
		a = 5;
		#100;
		a = 6;
		#100;
		a = 7;
		#100;
		a = 8;
		#100;
		a = 9;
		#100;
		a = 10;
		#100;
		a = 11;
		#100;
		a = 12;
		#100;
		a = 13;
		#100;
		a = 14;
		#100;
		a = 15;
		#100;
	end
endmodule
