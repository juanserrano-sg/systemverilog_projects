
/******************************************************************
* Description
*
* I2C Master Generator
*
* Author: Juan Antonio Serrano Gomez
* email : antonio.serrano@cinvestav.mx
* Date  :	09/06/2023
******************************************************************/


module I2C_GEN(
	input clk,
	inout SDA,
	output SCL
	
);
	
	logic [7:0] dataRx;				// Sores the data received from the slave
	int i;
	logic SDA_INT = 1'b1;			// SDA internal signal
	logic SCL_INT = 1'b1;			// SCL internal signal
	logic [3:0] cnt = 0;			// Clock (clk) TICs counter
	logic [3:0] bitCnt = 0;			// Used to counts the bits transmitted/received to/from the slave
	logic wr = 1'b0; 				// Asserted when DATA is trasmitted to the slave 
	logic rd = 1'b0;    			// Asserted when DATA is received from the slave
	localparam TICS = 5;
	
	assign SCL = SCL_INT;           
	assign SDA = !(SDA_INT) ? 1'b0 : 1'bz;
	
	// This task is used to generate the START pulse
	task start;  	
		begin
		    SCL_INT = 1'b1;
			SDA_INT = 1'b1;
			for (i=0; i<3; i++) begin
				cnt = 0;
				while (cnt < TICS) begin
					@(posedge clk)
					cnt++;
				end
				if (!wr && !rd) begin	// START pulse generation 
					i = 3;
					SDA_INT = 1'b0;
				end
				else if (wr) begin		// START pulse generation after data transmitted to the slave
					SCL_INT = ~SCL_INT;
					if (i == 2) begin
						SDA_INT = 1'b0;
						i = 3;
					end
				end
			    else if (rd) begin		// START pulse generation after data received from the slave
					SDA_INT = 1'b0;				
					i = 3;
				end					
			end
			wr = 1'b0;
			rd = 1'b0;
		end
	endtask
	
	// This task is used to generate the STOP pulse
	task stop; 
		begin
		    SCL_INT = 1'b1;
			SDA_INT = 1'b0;
			for (i=0; i<3; i++) begin
				cnt = 0;
				while (cnt < TICS) begin	
					@(posedge clk)
					cnt++;
				end
				if (!wr && !rd) begin	 	// STOP pulse generation 
					SDA_INT = 1'b1;                 
					i =3;               
				end                         
				else if (wr) begin		  	// STOP pulse generation after data transmitted to the slave  
					SCL_INT = ~SCL_INT;     
					if (i == 2) begin  
						SDA_INT = 1'b1;  
						SCL_INT = 1'b1;           
					end
				end
				else if (rd) begin			// STOP pulse generation after data received from the slave
					SDA_INT = 1'b1; 
					i = 3;
				end
			end
			wr = 1'b0;
			rd = 1'b0;
		end
	endtask
	
	// This task is used to transmit data to the slave
	task txData;
		input [7:0] data ;
		begin
			wr = 1'b1;
			cnt = 0;
			bitCnt = 8;
			SCL_INT = 1'b1;
			while (bitCnt > 0 || !SCL_INT) begin // Wait until 8 bit are transmitted to the slave
				while (cnt < TICS) begin
					@(posedge clk)
					cnt++;
				end
				
				cnt = 0;
				SCL_INT = ~SCL_INT;
				if (!SCL_INT) begin			 
				    bitCnt--;
					SDA_INT = data[bitCnt];	  	// One bit is transmitted to the slave
					
				end
			end	
			cnt = 0;
			while (cnt < TICS) begin     		    
				@(posedge clk)
				cnt++;
			end
			SDA_INT = 1'b1;  							
			SCL_INT = 1'b0;						// ACK bit is generated by the slave
			cnt = 0;
			while (cnt < TICS) begin         
				@(posedge clk)
				cnt++;
			end
			SCL_INT = 1'b1;						// ACK bit is read
			if (SDA) 	
				$display("NACK received");			
		end
	endtask
	
	// This task is used to receive data from the slave
	task rxData; input [7:0] dataExp;
		begin
			rd = 1'b1;
			cnt = 0;
			bitCnt = 8;
			SCL_INT = 1'b1;
			while (bitCnt > 0) begin 					// Wait until 8 bit are received from the slave
				while (cnt < TICS) begin
					@(posedge clk)
					cnt++;
				end
				cnt = 0;
				SCL_INT = ~SCL_INT;
				if (SCL_INT) begin	
					bitCnt--;			    
					dataRx[bitCnt] = SDA;				// One bit is received from the slave					
				end
			end	
			if (dataRx != dataExp)
				$display("ERROR at time %g: Expected data (%h) does not match Read data (%h)", $time, dataExp, dataRx);
				
			cnt = 0;	
			while (cnt < TICS) begin					
				@(posedge clk)
				cnt++;
			end
			SCL_INT = 1'b0;								
			SDA_INT = 1'b0;								// ACK bit is generated to the slave
			cnt = 0;	
			while (cnt < TICS) begin
				@(posedge clk)
				cnt++;
			end
			SCL_INT = 1'b1;								// ACK bit is read by the slave
		end
	endtask
	
endmodule
